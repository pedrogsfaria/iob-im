   // IM
   input [9:0] 	   im_pixel_x,
   input [9:0] 	   im_pixel_y,	
   output [11:0]   im_rgb,
