   // IM
   input [9:0] 	   pixel_x,
   input [9:0] 	   pixel_y,	
   output [11:0]   rgb,
